`timescale 1 ns / 1 ps

`include "transaction.sv"
`include "generator.sv"
`include "Driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "pico_intf.sv"
`include "env.sv"
`include "test_layered.sv"
`include "test_top.sv"
`include "picorv32.v"