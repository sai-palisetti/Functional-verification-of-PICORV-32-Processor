class insr_cover 


function new( );
   
  endfunction


covergroup cg;
	opcode	:	coverpoint mem

endgroup

endclass